library ieee;
USE ieee.numeric_std.all;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
--use std.textio.all; --  Imports the standard textio package.


--  A testbench has no ports.
   entity sum_data_chk_tb is
   end sum_data_chk_tb;
     
   architecture behav of sum_data_chk_tb is
      --  Declaration of the component that will be instantiated.
      component sum_data_chk
         port(
            Grs         : in std_logic;
            sum_in      : in std_logic_vector(63 downto 0);
            chan        : in std_logic_vector(5 downto 0);
            stat_msec   : in std_logic_vector(6 downto 0);
            prn_run     : in std_logic;
            stat_start  : in std_logic;
            OneMsec     : in std_logic;
            C125        : in std_logic;
            ecnt        : out std_logic_vector(7 downto 0);
            stat_p3     : out std_logic_vector(23 downto 0);
            stat_p1     : out std_logic_vector(23 downto 0);
            stat_m1     : out std_logic_vector(23 downto 0);
            stat_m3     : out std_logic_vector(23 downto 0);
            stat_rdy    : out std_logic
           );
      end component;

        --  Specifies which entity is bound with the component.
       for sum_data_chk_0: sum_data_chk use entity work.sum_data_chk;

        signal Grs_sig        : std_logic;
        signal sum_in_sig     : std_logic_vector(63 downto 0);
        signal chan_sig       : std_logic_vector(5 downto 0);
        signal stat_msec_sig  : std_logic_vector(6 downto 0);
        signal prn_run_sig    : std_logic;
        signal stat_start_sig : std_logic;
        signal OneMsec_sig    : std_logic;
        signal C125_sig       : std_logic;
        signal ecnt_sig       : std_logic_vector(7 downto 0);
        signal stat_p3_sig    : std_logic_vector(23 downto 0);
        signal stat_p1_sig    : std_logic_vector(23 downto 0);
        signal stat_m1_sig    : std_logic_vector(23 downto 0);
        signal stat_m3_sig    : std_logic_vector(23 downto 0);
        signal stat_rdy_sig   : std_logic;

     begin
        --  Component instantiation.
       sum_data_chk_0: sum_data_chk
          port map (
            Grs        => Grs_sig,
            sum_in     => sum_in_sig,
            chan       => chan_sig,
            stat_msec  => stat_msec_sig,
            prn_run    => prn_run_sig,
            stat_start => stat_start_sig,
            OneMsec    => OneMsec_sig,
            C125       => C125_sig,
            ecnt       => ecnt_sig, 
            stat_p3    => stat_p3_sig,
            stat_p1    => stat_p1_sig,
            stat_m1    => stat_m1_sig,
            stat_m3    => stat_m3_sig,
            stat_rdy   => stat_rdy_sig
         );
     
        --  This process does the real job.
        process
--           variable s : line;

           type pattern_type is record
              --  The inputs and outputs of the circuit
              sum_in     : std_logic_vector(63 downto 0);
              chan       : std_logic_vector(5 downto 0);
              stat_msec  : std_logic_vector(6 downto 0);
              prn_run    : std_logic;
              stat_start : std_logic;
              OneMsec    : std_logic;
              C125       : std_logic;
              ecnt       : std_logic_vector(7 downto 0);
              stat_p3    : std_logic_vector(23 downto 0);
              stat_p1    : std_logic_vector(23 downto 0);
              stat_m1    : std_logic_vector(23 downto 0);
              stat_m3    : std_logic_vector(23 downto 0);
              stat_rdy   : std_logic;
           end record;
           --  The patterns to apply.
           type pattern_array is array (natural range <>) of pattern_type;
           constant patterns : pattern_array :=
             --sum_in              chan     stat_msec prn_run
                                                            --stat_start
                                                                --OneMsec
                                                                    --C125
                                                                       --ecnt      stat_p3                    stat_p1                  stat_m1                   stat_m3                     stat_rdy
              --check 32:2 mux
             ((X"0000000000000001","000000","0000001",'0', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --1 ns
              (X"0000000000000001","000000","0000001",'0', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --2 ns
              (X"0000000000000008","000010","0000001",'0', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --3 ns
              (X"0000000000000008","000010","0000001",'0', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --4 ns
              (X"0000000000000010","000100","0000001",'0', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --5 ns
              (X"0000000000000010","000100","0000001",'0', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --6 ns
              (X"0000000000000080","000110","0000001",'0', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --7 ns
              (X"0000000000000080","000110","0000001",'0', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --8 ns
              (X"0000000000000100","001000","0000001",'0', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --9 ns
              (X"0000000000000100","001000","0000001",'0', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --10 ns
              (X"0000000000000800","001010","0000001",'0', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --11 ns
              (X"0000000000000800","001010","0000001",'0', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --12 ns
              (X"0000000000001000","001100","0000001",'0', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --13 ns
              (X"0000000000001000","001100","0000001",'0', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --14 ns
              (X"0000000000002000","001100","0000001",'0', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --15 ns
              (X"0000000000002000","001100","0000001",'0', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --16 ns
              (X"4000000000000000","111110","0000001",'0', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --17 ns
              (X"4000000000000000","111110","0000001",'0', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --18 ns
              (X"C000000000000000","111110","0000001",'0', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --19 ns
              (X"C000000000000000","111110","0000001",'0', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --20 ns
              (X"4000000000000000","111110","0000001",'0', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --21 ns
              (X"4000000000000000","111110","0000001",'0', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --22 ns
              --test 2:1 mux
              (X"8000000000000000","111111","0000001",'0', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --23 ns
              (X"8000000000000000","111111","0000001",'0', '1','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --24 ns
              (X"8000000000000000","111110","0000001",'0', '1','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --25 ns
              (X"8000000000000000","111110","0000001",'0', '1','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --26 ns
              (X"4000000000000000","111111","0000001",'0', '1','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --27 ns
              (X"4000000000000000","111111","0000001",'0', '1','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --28 ns
              --test prg; prn_run <= '1'
              (X"4000000000000000","111110","0000001",'1', '1','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --29ns
              (X"4000000000000000","111110","0000001",'1', '1','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --30ns
              (X"4000000000000000","111110","0000001",'1', '1','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --31ns             
              (X"4000000000000000","111110","0000001",'1', '1','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --32ns             
                  --initialize: pulse OneMsec
              (X"4000000000000000","111110","0000001",'1', '1','1','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --33ns            
              (X"4000000000000000","111110","0000001",'1', '1','1','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --34ns             
                  -- load prg; takes 35 clocks
              (X"4000000000000000","111110","0000001",'1', '1','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '1'),  --35ns
              (X"4000000000000000","111110","0000001",'1', '1','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --36ns
              (X"4000000000000000","111110","0000001",'1', '1','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --37ns
              (X"4000000000000000","111110","0000001",'1', '1','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --38ns
              (X"4000000000000000","111110","0000001",'1', '1','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --39ns
              (X"4000000000000000","111110","0000001",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --40ns
              (X"4000000000000000","111110","0000001",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --41ns
              (X"4000000000000000","111110","0000001",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --42ns
              (X"4000000000000000","111110","0000001",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --43ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --45ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --46ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --47ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --48ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --47ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --48ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --49ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --50ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --51ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --52ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --53ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --54ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --55ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --56ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --57ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --58ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --59ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --60ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --61ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --62ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --63ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --64ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --65ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --66ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --67ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --68ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --69ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --70ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --71ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --72ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --73ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --74ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --75ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --76ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --77ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --78ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --79ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --80ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --81ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --82ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --83ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --84ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --85ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --86ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --87ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --88ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --89ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --90ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --91ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --92ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --93ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --94ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --95ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --96ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --97ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --98ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --99ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --100ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --101ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --102ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --103ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --104ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --105ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --106ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --107ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --108ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --109ns
              --test error counter; should count up except for one clock; i.e., stuck at count = 2 for 2 counts, otherwise increments
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --110ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --111ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --112ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --113ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --114ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --115ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --116ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --117ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --118ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --119ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --120ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --121ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --122ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --123ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --124ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --125ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --126ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --127ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --128ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --129ns
              --latch count and start PRN initialization again
              (X"4000000000000000","111110","0000011",'1', '0','1','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --130ns
              (X"4000000000000000","111110","0000011",'1', '0','1','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --131ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --132ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --133ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --134ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --135ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --136ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --137ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --138ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --139ns
              --let PRG initialize and this time and then insert a string of zeros so we can watch the zero counter operate
              -- set to 4 so we can see something in a finite amount of time
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --140ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --141ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --142ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --143ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --144ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --145ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --146ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --147ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --148ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --149ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --150ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --151ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --152ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --153ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --154ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --155ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --156ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --157ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --158ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --159ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --160ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --161ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --162ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --163ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --164ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --165ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --166ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --167ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --168ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --169ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --170ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --171ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --172ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --173ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --174ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --175ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --176ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --177ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --178ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --179ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --180ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --181ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --182ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --183ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --184ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --185ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --186ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --187ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --188ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --189ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --190ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --191ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --192ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --193ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --194ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --195ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --196ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --149ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --197ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --198ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --199ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --200ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --201ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --202ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --203ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --204ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --205ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --206ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --207ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --208ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --209ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --210ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --211ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --212ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --213ns
              (X"4000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --214ns
              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --215ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --216ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --217ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --218ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --219ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --220ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --221ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --222ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --223ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --224ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --225ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --226ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --227ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --228ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --229ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --230ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --231ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --232ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --233ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --234ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --235ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --236ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --237ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --238ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --239ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --240ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --241ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --242ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --243ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --244ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --245ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --246ns
              (X"8000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --247ns
              (X"8000000000000000","111110","0000011",'1', '0','0','1',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0'),  --248ns

              (X"4000000000000000","111110","0000011",'1', '0','0','0',"00000000", "000000000000000000000001", "000000000000000000000001","000000000000000000000001","000000000000000000000001", '0')   --249ns
             );
        begin
--           write (s, String'("at begin in test process"));
--           writeline (output, s);
--WAIT FOR 100 ns;

--just to get started
   C125_sig    <= '0';
   Grs_sig     <= '0';
   wait for 1 ns;
   Grs_sig     <= '1';
   wait for 1 ns;
   C125_sig    <= '1';
   wait for 1 ns;
   Grs_sig     <= '0';
   wait for 1 ns;
   C125_sig    <= '0';
--init_sig    <= '0';
--td_mode_sig <= "010";

--           write (s, String'("after initialization in test process"));
--           writeline (output, s);
--report "msg 3";
--wait for 1 ms;
--report "msg 4";
--           write (s, String'("Start of Test Data Generator Test Bench"));
--           writeline (output, s);

           --  Check each pattern.
           for i in patterns'range loop
              --  Set the inputs.
              C125_sig       <= patterns(i).C125;
              chan_sig       <= patterns(i).chan;
              stat_start_sig <= patterns(i).stat_start;
              OneMsec_sig    <= patterns(i).OneMsec;
              sum_in_sig     <= patterns(i).sum_in;
              prn_run_sig    <= patterns(i).prn_run;
              stat_start_sig <= patterns(i).stat_start;
              stat_msec_sig  <= patterns(i).stat_msec;
--           write (s, String'("msg2"));
--           writeline (output, s);
              wait for 1 ns;
--           write (s, String'("msg3"));
--           writeline (output, s);

              --  Check the outputs.

--              assert ecnt_sig = patterns(i).ecnt
--                 report "bad prg value" severity error;

           end loop;
--           write (s, String'("End first test loop"));
--           writeline (output, s);

          --for i in 0 to 3000000 loop
          --    wait for 1 ns;
          --    clk_sig  <= '1';
          --    wait for 1 ns;
          --    if (tst_data_sig = X"0000000000000001") then   
          --          write (s, String'("!!!!Found match!!!!"));
          --          writeline (output, s);
          --    end if;
          --    clk_sig  <= '0';
          -- end loop;

        --test the statistics logic
        wait for 10 ns;   --to get make an obvious place to start looking

        Grs_sig <= '1';   --initialize everything
        oneMsec_sig <= '0';
        C125_sig <= '0';
        wait for 1 ns;
        Grs_sig <= '0';

        wait for 1 ns;
        sum_in_sig    <= X"0000000000000002";    --set up to count minus threes for one msec
        chan_sig      <= "000000";
        stat_msec_sig <= "0000001";

        wait for 1 ns;   --start the sequence
        C125_sig       <= '0';
        stat_start_sig <= '1';

        wait for 1 ns;
        for i in 0 to 3 loop
           C125_sig       <= '0';
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
        end loop;

        C125_sig       <= '0';
        oneMsec_sig    <= '1';  --give a oneMsec pulse
        wait for 1 ns;   
        C125_sig       <= '1';
        oneMsec_sig    <= '1';
        wait for 1 ns;
        C125_sig       <= '0';
        oneMsec_sig    <= '0';  --give a oneMsec pulse
        wait for 1 ns;   
        C125_sig       <= '1';
        oneMsec_sig    <= '0';
        wait for 1 ns;
        
        for i in 0 to 21 loop   --count for 21 clocks
           C125_sig       <= '0';
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
        end loop;

        C125_sig       <= '0';
        oneMsec_sig    <= '1';  --give a oneMsec pulse
        wait for 1 ns;   
        C125_sig       <= '1';
        oneMsec_sig    <= '1';
        wait for 1 ns;
        C125_sig       <= '0';
        oneMsec_sig    <= '0'; 
        wait for 1 ns;   
        C125_sig       <= '1';
        oneMsec_sig    <= '0';
        wait for 1 ns;

        for i in 0 to 3 loop     --give a couple more clocks
           C125_sig       <= '0';
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
        end loop;

        --bigger test: should result in 1:2:3:4 ratio of counts, except for starting offset
        wait for 1 ns;          --bring stat_start low and then high
        C125_sig       <= '0';
        stat_start_sig <= '0';
        wait for 1 ns;
        C125_sig       <= '1';
        wait for 1 ns;
        C125_sig       <= '0';
        stat_start_sig <= '1';
        wait for 1 ns;
        C125_sig       <= '1';
        wait for 1 ns;
        C125_sig       <= '0';

        wait for 1 ns;          --give a few clocks
        for i in 0 to 3 loop
           C125_sig       <= '0';
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
        end loop;


        C125_sig       <= '0';   --give a oneMsec pulse to start the counting
        oneMsec_sig    <= '1';  
        wait for 1 ns;   
        C125_sig       <= '1';
        oneMsec_sig    <= '1';
        wait for 1 ns;
        C125_sig       <= '0';
        oneMsec_sig    <= '0'; 
        wait for 1 ns;   
        C125_sig       <= '1';
        oneMsec_sig    <= '0';
        wait for 1 ns;

        for i in 0 to 5 loop       --bigger loop to generate ratio of counts
           sum_in_sig    <= X"0000000000000002";     --minus 3      
           C125_sig       <= '0';                    --one clock
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           sum_in_sig    <= X"0000000000000003";     --minus 1      
           C125_sig       <= '0';                    --two clocks
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           C125_sig       <= '0';                   
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           sum_in_sig    <= X"0000000000000000";     --plus 1      
           C125_sig       <= '0';                    --three clocks
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           C125_sig       <= '0';                   
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           C125_sig       <= '0';                   
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           sum_in_sig    <= X"0000000000000001";     --plus 3      
           C125_sig       <= '0';                    --four clocks
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           C125_sig       <= '0';                   
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           C125_sig       <= '0';                   
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           C125_sig       <= '0';                   
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;      
        end loop;

        C125_sig       <= '0';   --give a oneMsec pulse to end the counting
        oneMsec_sig    <= '1';  
        wait for 1 ns;   
        C125_sig       <= '1';
        oneMsec_sig    <= '1';
        wait for 1 ns;
        C125_sig       <= '0';
        oneMsec_sig    <= '0'; 
        wait for 1 ns;   
        C125_sig       <= '1';
        oneMsec_sig    <= '0';
        wait for 1 ns;

        wait for 1 ns;          --give a few clocks
        for i in 0 to 3 loop
           C125_sig       <= '0';
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
        end loop;


        --even bigger test: should result in 1:2:3:4 ratio of counts, except for starting offset
        -- plus should count for 3 msec
        wait for 1 ns;          --bring stat_start low and then high
        C125_sig       <= '0';
        stat_start_sig <= '0';
        stat_msec_sig  <= "0000011"; --3 msec request

        wait for 1 ns;
        C125_sig       <= '1';
        wait for 1 ns;
        C125_sig       <= '0';
        stat_start_sig <= '1';
        wait for 1 ns;
        C125_sig       <= '1';
        wait for 1 ns;
        C125_sig       <= '0';

        wait for 1 ns;          --give a few clocks
        for i in 0 to 3 loop
           C125_sig       <= '0';
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
        end loop;

        outer: for j in 0 to 4 loop

        C125_sig       <= '0';   --give a oneMsec pulse to start the counting
        oneMsec_sig    <= '1';   --note that this results in 2 extra +3 counts 
        wait for 1 ns;   
        C125_sig       <= '1';
        oneMsec_sig    <= '1';
        wait for 1 ns;
        C125_sig       <= '0';
        oneMsec_sig    <= '0'; 
        wait for 1 ns;   
        C125_sig       <= '1';
        oneMsec_sig    <= '0';
        wait for 1 ns;

        inner: for i in 0 to 5 loop       --loop to generate ratio of counts
           sum_in_sig    <= X"0000000000000002";     --minus 3      
           C125_sig       <= '0';                    --one clock
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           sum_in_sig    <= X"0000000000000003";     --minus 1      
           C125_sig       <= '0';                    --two clocks
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           C125_sig       <= '0';                   
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           sum_in_sig    <= X"0000000000000000";     --plus 1      
           C125_sig       <= '0';                    --three clocks
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           C125_sig       <= '0';                   
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           C125_sig       <= '0';                   
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           sum_in_sig    <= X"0000000000000001";     --plus 3      
           C125_sig       <= '0';                    --four clocks
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           C125_sig       <= '0';                   
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           C125_sig       <= '0';                   
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
           C125_sig       <= '0';                   
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;      
        end loop inner;
      end loop outer;

        wait for 1 ns;          --give a few clocks
        for i in 0 to 3 loop
           C125_sig       <= '0';
           wait for 1 ns;
           c125_sig       <= '1';
           wait for 1 ns;
        end loop;

        
        


           assert false report "end of test" severity note;
           --  Wait forever; this will finish the simulation.
           wait;


        end process;
     end behav;
