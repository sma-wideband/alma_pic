-------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;
-------------------------------------------------------

--This entity packs the sum data according to the number of channels to be recorded
--See the ICD with computing for cool graphics showing the details and comments in the
--code below for additional details

entity header_collator is
 port(
	 -- timing reference signals 
	 C125        : in std_logic; 	
	 TE			 : in std_logic; 	
		
   --data from which to form header
     --packet serial number from data_write_ctrl
     PSN         : in std_logic_vector(63 downto 0); 

     --bad frame indicator bit from microprocessor
     badFrame    : in std_logic; 

     --time info from timing generator
     SFRE        : in std_logic_vector(29 downto 0); --seconds from ref. epoch
     FrameNum    : in std_logic_vector(23 downto 0); --data frame number

     --data from microprocessor interface
     refEpoch : in std_logic_vector(5 downto 0);
     nchan : in std_logic_vector(4 downto 0);
     frameLength : in std_logic_vector(23 downto 0);
     threadID    : in std_logic_vector(9 downto 0);
     stationID   : in std_logic_vector(15 downto 0);
     magicWord   : in std_logic_vector(23 downto 0);
     statusWord  : in std_logic_vector(31 downto 0); 
      
   --data output of collator to header_fifo
     coll_out    : out std_logic_vector(63 downto 0);

   --control of the header mux from data_write_control
     hdr_sel     : in std_logic_vector(2 downto 0);
	 
   --data output of collator to C167
     coll_out_c167    : out std_logic_vector(7 downto 0);   
   --control of the header mux from C167
     hdr_sel_c167     : in std_logic_vector(5 downto 0)   
	 
	 
);
end header_collator;

architecture arch of header_collator is
  --signal definitions
    --the output of the collator
      signal coll_out_sig: std_logic_vector(63 downto 0) := X"1000_2000_3000_0001";
	  signal coll_out_c167_sig: std_logic_vector(7 downto 0) := X"00";
      
    --the header words that are comprised of multiple quantities, as defined in the VDIF packet definition
      signal word0      : std_logic_vector(31 downto 0):= X"4000_0000";
      signal word1      : std_logic_vector(31 downto 0):= X"5000_0000";
      signal word2      : std_logic_vector(31 downto 0):= X"6000_0000";
      signal word3      : std_logic_vector(31 downto 0):= X"7000_0000";
      signal word4      : std_logic_vector(31 downto 0):= X"8000_0000";
      
      --long (64-bit) words comprised of pairs of the above words for sending to fifo
      signal lWord0      : std_logic_vector(63 downto 0);
      signal lWord1      : std_logic_vector(63 downto 0);
      signal lWord2      : std_logic_vector(63 downto 0);
      signal lWord3      : std_logic_vector(63 downto 0);
      signal lWord4      : std_logic_vector(63 downto 0);  

	  signal lWord0_register      : std_logic_vector(63 downto 0);
	  signal lWord1_register      : std_logic_vector(63 downto 0);
	  signal lWord2_register      : std_logic_vector(63 downto 0);
	  signal lWord3_register      : std_logic_vector(63 downto 0);
	  signal lWord4_register      : std_logic_vector(63 downto 0);
	  
	  signal TE_s		 : std_logic;

  begin
    --output of mux
    coll_out <= coll_out_sig;
	coll_out_c167 <= coll_out_c167_sig;
  
    --form 32-bit words from various pieces of info
    word0    <= badFrame & '0' & SFRE;
    word1    <= "00" & refEpoch & FrameNum;
    word2    <= "000" & nchan & frameLength;
    word3    <= "000001" & threadID & stationID;
    word4    <= X"02" & magicWord;
    --word5    <= statusWord;
    --word 6 and 7 are a repeat of the PSN
    
    --form 64-bit words from 32-bit words
    lWord0   <= PSN(31 downto 0) & PSN(63 downto 32);    
    lWord1   <= word0 & word1;
    lWord2   <= word2 & word3;
    lWord3   <= word4 & statusWord;
    lWord4   <= PSN(31 downto 0) & PSN(63 downto 32);    
    
    mux: process(Hdr_sel, lWord0, lWord1, lWord2, lWord3, lWord4)
    begin
        case Hdr_sel is                 -- data selection signals
      	  when "000"  => coll_out_sig <= lWord0;
        	when "001"  => coll_out_sig <= lWord1;     
        	when "010"  => coll_out_sig <= lWord2;
        	when "011"  => coll_out_sig <= lWord3;
        	when "100"  => coll_out_sig <= lWord4;
        	when others => coll_out_sig <= X"0000_0000_0000_0000";
       end case;
    end process;
	
	
	process(C125,TE)
	begin
		if c125='1' and c125'event then			
			TE_s <= TE; 
		end if;
    end process;	
	
	
	capture_upon_te_rising_edge: process(C125,TE,TE_s,lWord0,lWord1,lWord2,lWord3,lWord4)
	begin
		if c125='1' and c125'event then			
			if TE='1' and TE_s='0' then
				lWord0_register <= lWord0;
				lWord1_register <= lWord1;
				lWord2_register <= lWord2;
				lWord3_register <= lWord3;
				lWord4_register <= lWord4;
			 end if;	
		end if;				
	end process;
	
	mux_c167: process(Hdr_sel_c167,lWord0,lWord1,lWord2,lWord3,lWord4)
	begin
		case Hdr_sel_c167 is
			when "000000" => coll_out_c167_sig <= lWord0_register(7 downto 0);		-- 0
			when "000001" => coll_out_c167_sig <= lWord0_register(15 downto 8);		-- 1
			when "000010" => coll_out_c167_sig <= lWord0_register(23 downto 16);	-- 2
			when "000011" => coll_out_c167_sig <= lWord0_register(31 downto 24);	-- 3
			when "000100" => coll_out_c167_sig <= lWord0_register(39 downto 32);	-- 4
			when "000101" => coll_out_c167_sig <= lWord0_register(47 downto 40);	-- 5
			when "000110" => coll_out_c167_sig <= lWord0_register(55 downto 48);	-- 6
			when "000111" => coll_out_c167_sig <= lWord0_register(63 downto 56);	-- 7
			when "001000" => coll_out_c167_sig <= lWord1_register(7 downto 0);		-- 0
			when "001001" => coll_out_c167_sig <= lWord1_register(15 downto 8);		-- 1
			when "001010" => coll_out_c167_sig <= lWord1_register(23 downto 16);	-- 2
			when "001011" => coll_out_c167_sig <= lWord1_register(31 downto 24);	-- 3
			when "001100" => coll_out_c167_sig <= lWord1_register(39 downto 32);	-- 4
			when "001101" => coll_out_c167_sig <= lWord1_register(47 downto 40);	-- 5
			when "001110" => coll_out_c167_sig <= lWord1_register(55 downto 48);	-- 6
			when "001111" => coll_out_c167_sig <= lWord1_register(63 downto 56);	-- 7			
			when "010000" => coll_out_c167_sig <= lWord2_register(7 downto 0);		-- 0
			when "010001" => coll_out_c167_sig <= lWord2_register(15 downto 8);		-- 1
			when "010010" => coll_out_c167_sig <= lWord2_register(23 downto 16);	-- 2
			when "010011" => coll_out_c167_sig <= lWord2_register(31 downto 24);	-- 3
			when "010100" => coll_out_c167_sig <= lWord2_register(39 downto 32);	-- 4
			when "010101" => coll_out_c167_sig <= lWord2_register(47 downto 40);	-- 5
			when "010110" => coll_out_c167_sig <= lWord2_register(55 downto 48);	-- 6
			when "010111" => coll_out_c167_sig <= lWord2_register(63 downto 56);	-- 7
			when "011000" => coll_out_c167_sig <= lWord3_register(7 downto 0);		-- 0
			when "011001" => coll_out_c167_sig <= lWord3_register(15 downto 8);		-- 1
			when "011010" => coll_out_c167_sig <= lWord3_register(23 downto 16);	-- 2
			when "011011" => coll_out_c167_sig <= lWord3_register(31 downto 24);	-- 3
			when "011100" => coll_out_c167_sig <= lWord3_register(39 downto 32);	-- 4
			when "011101" => coll_out_c167_sig <= lWord3_register(47 downto 40);	-- 5
			when "011110" => coll_out_c167_sig <= lWord3_register(55 downto 48);	-- 6
			when "011111" => coll_out_c167_sig <= lWord3_register(63 downto 56);	-- 7			
			when "100000" => coll_out_c167_sig <= lWord4_register(7 downto 0);		-- 0
			when "100001" => coll_out_c167_sig <= lWord4_register(15 downto 8);		-- 1
			when "100010" => coll_out_c167_sig <= lWord4_register(23 downto 16);	-- 2
			when "100011" => coll_out_c167_sig <= lWord4_register(31 downto 24);	-- 3
			when "100100" => coll_out_c167_sig <= lWord4_register(39 downto 32);	-- 4
			when "100101" => coll_out_c167_sig <= lWord4_register(47 downto 40);	-- 5
			when "100110" => coll_out_c167_sig <= lWord4_register(55 downto 48);	-- 6
			when "100111" => coll_out_c167_sig <= lWord4_register(63 downto 56);	-- 7
			when others => coll_out_c167_sig   <= X"00";
		end case;	
	end process;

  end arch;

      
   
